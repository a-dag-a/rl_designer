* Common Source Amplifier

* Define parameters
.param param__VDD = 12V
.param param__VSS = 0V
.param param__VGS = 2.5V
.param param__RD = 2k
.param param__RS = 1k
.param param__RL = 10k
.param param__C1 = 10u
.param param__C2 = 10u
.param param__gm = 2e-3
.param param__ro = 100k

* Voltage sources
VDD vdd 0 DC {param__VDD}
VSS 0 vss DC {param__VSS}
VGS gate 0 DC {param__VGS}

* Input source
Vin in 0 AC 1

* Transistor model
.model NMOS NMOS(VTO=1 KP=1e-4)

* NMOS transistor
M1 drain gate source 0 NMOS

* Resistors and capacitors
RD drain vdd {param__RD}
RS source vss {param__RS}
RL drain out {param__RL}
C1 in gate {param__C1}
C2 out vss {param__C2}

* Load resistor
Rload out 0 1Meg

* AC analysis
.ac dec 10 1 1Meg

* Print AC analysis results
.print ac v(out)

.end
